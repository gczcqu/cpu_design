`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2017/11/07 10:58:03
// Design Name: 
// Module Name: mips
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module mips(
	input wire clk,rst,
	output wire[31:0] pcF,
	input wire[31:0] instrF,
	output wire memwriteM,
	output wire[31:0] data_addr,writedataM,
	input wire[31:0] readdataM,
	output wire [3:0]data_wenM
    );
	
	wire [5:0] opD,functD;
	wire regdstE,alusrcE,pcsrcD,signimmnextD,memtoregE,hiloregwriteE,hiloregreadE,memtoregM,memtoregW,
			regwriteE,regwriteM,regwriteW,hiloregreadW;
	wire [4:0] alucontrolE;
	wire flushE,equalD;
	wire [2:0]l_s_typeM;
	controller c(
		clk,rst,
		//decode stage
		opD,functD,
		pcsrcD,branchD,equalD,jumpD,
		
		//execute stage
		flushE,
		memtoregE,alusrcE,
		regdstE,regwriteE,	
		alucontrolE,
		hiloregwriteE,
		hiloregreadE,
		hiloregreadW,
		signimmnextD,
		//mem stage
		memtoregM,memwriteM,
		regwriteM,
		l_s_typeM,
		//write back stage
		memtoregW,regwriteW
		);
	datapath dp(
		clk,rst,
		//fetch stage
		pcF,
		instrF,
		//decode stage
		pcsrcD,branchD,
		jumpD,
		equalD,
		opD,functD,
		//execute stage
		memtoregE,
		alusrcE,regdstE,
		regwriteE,
		alucontrolE,
		hiloregwriteE,
		hiloregreadE,
		hiloregreadW,
		signimmnextD,
		flushE,
		//mem stage
		memtoregM,
		regwriteM,
		data_addr,writedataM,data_wenM,
		readdataM,
		l_s_typeM,
		//writeback stage
		memtoregW,
		regwriteW
	    );
	
endmodule
